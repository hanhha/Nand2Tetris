// HMTH (c)
// Instruction fetch - Instruction decode

module IfId (
);
endmodule
// EOF
