// HMTH (c)
// Memory Access - Read data

module Mr (
);
endmodule
// EOF
