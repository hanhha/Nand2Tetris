// HMTH (c)
// Memory Access

module Ma (
);
endmodule
// EOF
