// HMTH (c)
// Memory Access - Write data

module Mw (
);
endmodule
// EOF
